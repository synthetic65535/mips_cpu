parameter OP_R = 6'b000000;
parameter OP_ADDI = 6'b001000;
parameter OP_BEQ = 6'b000100;
parameter OP_BNE = 6'b000101;
parameter OP_LW = 6'b100011;
parameter OP_SW = 6'b101011;

parameter OPR_NOP = 6'b000000;
parameter OPR_ADD = 6'b100000;
parameter OPR_SUB = 6'b100010;

parameter ALU_ADD = 8'd00;
parameter ALU_SUB = 8'd01;

parameter R00 = 5'd00;
parameter R01 = 5'd01;
parameter R02 = 5'd02;
parameter R03 = 5'd03;
parameter R04 = 5'd04;
parameter R05 = 5'd05;
parameter R06 = 5'd06;
parameter R07 = 5'd07;
parameter R08 = 5'd08;
parameter R09 = 5'd09;
parameter R10 = 5'd10;
parameter R11 = 5'd11;
parameter R12 = 5'd12;
parameter R13 = 5'd13;
parameter R14 = 5'd14;
parameter R15 = 5'd15;
parameter R16 = 5'd16;
parameter R17 = 5'd17;
parameter R18 = 5'd18;
parameter R19 = 5'd19;
parameter R20 = 5'd20;
parameter R21 = 5'd21;
parameter R22 = 5'd22;
parameter R23 = 5'd23;
parameter R24 = 5'd24;
parameter R25 = 5'd25;
parameter R26 = 5'd26;
parameter R27 = 5'd27;
parameter R28 = 5'd28;
parameter R29 = 5'd29;
parameter R30 = 5'd30;
parameter R31 = 5'd31;
