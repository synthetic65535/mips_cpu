
module cpu (
  input [31:0] in,
  output reg [31:0] out,
  input load, clock
  );
  
  
  
endmodule
